-- --------------------------------------------------------------------
-- SPDX-License-Identifier: LGPL-3.0-or-later or CERN-OHL-W-2.0
-- prescaler.vhd is a part of Innervator.
-- --------------------------------------------------------------------







-- --------------------------------------------------------------------
-- END OF FILE: prescaler.vhd
-- --------------------------------------------------------------------