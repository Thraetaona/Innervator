-- NOTE: This was initially meant to be automated, but it was outright
-- impossible due to Vivado's noncompliance with the VHDL-2008 standard
-- for using allocators as to generate synth'able code.
-- See: network_parser.vhd

library ieee;
    use ieee.std_logic_1164.all; -- Added to fix ModelSim's errors

library config;
    context config.neural_context;


package network_params is
    -- NOTE: Use the boilerplate code in 'neural_typedefs.vhd' to bring
    -- attributes/groups to the constants (NOT unconstrained arrays)
    -- defined herein.
    constant NUM_NEURONS : integer_vector := (64, 20, 10);
    constant NUM_LAYERS  : natural := 2; -- Hidden & Output layers only

    -- Biases' 1-D arrays
    constant BIASES_1 : neural_array := 
        ("10110011","11101000","00111011","01011010","10111111","01100110","10010110","10101101","00011100","01101111","10001110","00010000","11011110","01111001","10010110","00000010","00100011","10010001","11011001","00010000");
    constant BIASES_2 : neural_array := 
        ("10011000","10010101","10111010","10101011","10011101","10100100","10011110","10011111","10100001","10011111");
    
    -- Weights' 1-D (NOT 2-D) array OF array (i.e., nested array)
    constant WEIGHTS_1 : neural_matrix := (
        ("00000111","11111110","00010000","00010011","00011001","00011010","00010101","00010000","11110101","11110011","00000000","00010000","00000010","11111001","00000011","11111011","00001101","11110010","00000100","00001000","11110111","11011101","11101100","00000010","11111101","00001111","00000100","00000000","11111000","00000011","11110010","00001100","11111101","11111001","00000111","00000100","00000010","00000001","00000011","00010000","11111101","11110100","11110010","11111111","11110000","00001101","00000110","00000101","00001010","11110101","00000001","00011001","00000000","11110010","00000100","00000100","11111101","11110010","00010100","00010011","11111000","11110011","00000101","00000100"),
        ("00001000","00000001","00000100","11110101","00000100","00001100","11110010","00001011","00000101","11110110","11110001","11111101","11110110","11110010","11111110","00001101","11110100","00000101","11110100","00000110","00001011","00000010","00001101","00001001","11111110","00000111","00001010","00000000","00001000","00000110","00001010","11110100","00000101","11110001","00001011","00000011","00000011","00000011","11110100","11110100","11110000","11111111","00001100","00001011","00010101","11111000","11111111","11110101","11111100","00001011","11111001","11110011","11110110","11111110","11110101","00001011","00000011","11111010","00000110","00001010","00001100","11110101","00000111","11111100"),
        ("00001000","11111001","00000101","00000110","00000000","11111100","11111110","11111111","11111001","00001100","00001000","11111010","00000010","11111101","00001101","11110010","00001011","11111001","00010110","00000001","00001110","11110001","11110110","00001000","11111101","11110111","00000010","11111011","11111101","11111000","11111001","11111010","11111010","00001010","00001001","00011101","00010011","11111111","00000000","11111110","00001110","00000011","00011101","00011000","00000011","00000001","11111001","00001000","00000010","00001100","00010001","00100010","00001010","00000111","00100000","00001101","00001001","00000001","11111110","11111111","00011010","00100111","00001101","11111011"),
        ("11111101","11110100","00001100","00000111","00010010","00010101","00000111","11111000","11110111","11110110","11110111","00001111","00000010","00010001","00001101","00001011","00000011","00000001","00000110","00001000","00100001","00001011","11111010","11110100","00001110","11110110","00010101","00100100","00011111","00001000","11111000","00000111","00001101","11111100","11111111","00010110","00100101","00001111","00000011","11111000","00000010","11110100","11111011","00000000","00010100","00010010","00000001","00000100","11111001","11110111","11111001","11110010","00001001","11111111","11101001","00000110","11110110","11111010","00001010","11111011","11111100","11101110","11111010","00000110"),
        ("00001111","00000101","00001010","11110110","00000100","00000100","00000111","11110110","00000111","00000111","00011111","00001011","00000110","11110101","00000010","00000011","11111111","00000101","00011000","00000001","11100100","00010101","00001000","00001100","00000010","00000100","00011000","00000101","00001001","00001010","00000101","00000001","11111001","00001110","00001100","11111100","11100110","11111001","00010100","00000001","00001101","00011000","00000111","11111111","00001100","00001001","00000011","11110011","00000101","11111001","00000000","11100001","00001001","11111011","11101000","00000110","11110001","00000011","00000101","00000011","00001101","11011100","11110111","11111111"),
        ("00000111","11110100","11110101","11111100","00001101","11110101","11110000","00001001","00000110","11111101","00000101","00001010","00000001","00001110","00001001","11111001","11111111","00000110","11111111","00000010","00001001","00010001","11111010","11111110","11111100","11111100","11111111","11111100","11111011","00001000","11110110","00000110","11110011","11111101","00001011","00001010","00010000","00001000","00001001","00001110","00001001","11111100","00010000","11110111","00001011","00000000","11111110","11111001","00000001","11111101","11110110","00000111","00000111","11111011","11110101","00000111","11111000","11111011","00001110","11111011","11111010","00001110","00001001","00000000"),
        ("11111100","00010001","00010101","00000110","00000101","00000100","00000100","11110100","11111011","00010001","00001011","00000010","11111010","00000001","00001011","11110011","11111011","00001110","00000100","00000000","11111100","11111001","00001010","00010000","00000011","00000011","11110011","00000000","00000111","11111010","00001101","00000100","11110000","00000101","00000000","00000111","00000111","00000001","11110010","11111111","00001110","00001011","11101111","00001000","11101111","11111110","00000101","11110010","00000001","00001000","00000000","00010011","00000100","11111100","00000101","00000001","00001000","00001111","00000001","00010000","00000100","00001101","00001010","11111110"),
        ("00000110","00000001","00001011","00001101","00000001","11110101","11110011","00000010","00000100","00000101","00001101","00001001","11111001","00000001","00010011","11111010","11110100","11110111","11111111","00000011","00001110","00011001","00011000","11110111","00001011","00000011","11111110","00000111","00011010","00010011","11111010","11111000","11110100","11111101","11101010","00001100","00000001","00001011","11110111","11111101","11111110","11111011","11110000","11101101","11101011","00000010","00010011","11111101","00000010","00001001","11111010","11111100","11110101","11111110","00001001","11110010","00001111","11111101","11110110","00000101","00000101","11111011","11111011","00001011"),
        ("11110001","11110000","00000100","11111011","11110001","11111011","00001010","00000010","11110010","11110100","11101110","11101111","00000110","11111000","11110011","11110111","00000011","00000011","11110111","00001010","00010110","00000111","00000101","00000010","00001111","00000101","00000101","11110110","00000000","00001001","00001101","00001111","00001101","11111000","00000101","11110001","00000110","00001000","11111000","00001011","11110001","00000111","11110000","00001110","00000110","11110100","00000011","11111010","11110111","11110011","11100011","00000110","00001011","11110100","11111010","11111011","00000001","00001001","11111001","00000101","00000011","11111000","11111100","11111101"),
        ("00000001","11111111","11101100","11111110","11110111","11101001","11101101","00000010","00000001","11110011","00000111","00000111","00001110","00001101","11110010","00001100","11110010","00000010","00001110","00011011","00000000","00000110","00001011","00000101","11111001","00000110","00000111","11110000","11110100","00001000","00001000","11110100","00001100","00001110","00001110","00010000","00010010","11101111","11111011","11111000","11110101","00000110","00100101","00011101","00001000","00000011","11110011","00000100","00001001","00000111","00001101","00010001","00011100","00011100","11111101","11110110","11110100","00000001","11110010","00010000","00011100","00001010","00011011","11111001"),
        ("00001111","00000111","00001110","00001001","00010000","00010101","00000000","00000001","11110010","00001000","11111111","00000010","00001000","00000100","11111001","11111001","11110101","11111110","11110101","11111110","00010001","00000111","00001001","11110001","00000010","11111110","11101101","00000000","00011000","11110101","11110100","11111100","11111100","11110110","11100101","00000100","00011000","11110110","11100101","11111100","11111100","11111011","11111100","00000001","00010111","11110001","00000000","00001000","11111000","00001000","00001011","00000001","00011100","00010110","00001111","11110111","11111010","00001110","00000001","11111110","00001110","00010001","00001110","00001110"),
        ("00000100","00001100","11111111","11111100","00001101","00000000","00001011","11110111","11110101","11111001","11111110","00001000","11111111","11111111","11110111","00000000","11111111","00000110","00000010","11111000","00000100","11111010","11110001","11111011","11110011","00000011","00000100","11110010","11110011","11111100","00001001","00001111","11110101","11110111","00001101","11111101","00001100","11110100","11110001","11110110","00001110","11111011","00000001","11110110","00001011","11111011","11110000","00000001","11110011","11111011","11110111","00000111","11110011","00001000","00000100","00000111","00000001","00001001","00000100","11111100","11111110","11110111","11110111","11110110"),
        ("11111000","11111011","00000000","00001000","00010001","00000100","11110101","11111101","00001011","11110111","00001001","11111001","11111111","11110101","00001001","00000011","11110111","00010010","00011010","11110111","00001000","00001111","11111100","00000111","00001011","11110001","00001101","00001011","11111100","11111010","11111110","00000001","00000001","11110001","11110011","11111011","11111000","11111110","00001010","00000101","00001010","11110001","11101001","11100101","00000001","00001010","11111000","00000110","00000101","00001001","11111001","11110100","11111011","11111010","11111011","11111101","11110001","11110101","00000110","00001011","00000000","00000101","00001001","11111101"),
        ("00000000","00001101","11110000","00000110","00001101","11110100","00001000","11111110","11111011","11111101","11111111","00001000","00010001","00000001","11111111","11111101","11111101","11111100","00001011","00001000","00000010","00010101","00010100","00000110","00000110","11111110","00010100","00000010","11111110","00011101","00011111","00001100","00000010","00001111","00001111","00001110","11110101","00101100","00011101","11110111","00000111","00000100","00001111","00011100","00010011","00000100","00011001","00000100","00000011","11111000","11111111","00001100","11110000","11110011","00001001","00000011","00001010","11111100","11111110","11111011","11100110","00000010","00000001","00000010"),
        ("11111001","11110011","00000000","00011100","00010011","00000110","00000011","00010000","00000110","11110011","00011001","00000111","00001010","00100001","00001000","00001001","11111110","00000111","11110110","11110010","11111001","00010100","00000011","00001110","11111001","11100000","11111000","11111010","11111000","00000100","00001000","00001000","11111000","11101101","00001011","00001101","00010101","00000100","11110111","11111100","00000010","00001001","00011101","11110001","11111100","00000011","00010100","00000100","11111000","00000000","00001100","00000010","11011111","00000011","00000110","00000110","11111011","11110010","11111000","00010011","00000110","11111110","11110000","00000001"),
        ("11110001","00001011","11110000","11110001","00000011","00000110","00000010","11110001","11111100","11111001","11101010","11111101","11101010","11111001","11111101","00001000","11111001","00000000","00100000","00010011","11110101","11101100","11110100","00010000","11110110","00001111","00010011","00100110","00010010","00000000","11110101","00001011","11110101","00000101","00001100","00010110","00000101","11111110","00000011","00000000","00000000","11111000","11110101","00000001","00011000","00000101","00000111","11110100","11110001","00000110","00001000","11101100","11100011","11110111","00000000","00001010","11111001","11110001","00000000","11110001","00000111","00000011","11110010","00000101"),
        ("00000100","11111111","00000110","11110011","11110110","00001001","11111111","11110111","11111001","11111110","00000011","11111111","11111000","11110001","00001001","00000111","00001010","11111001","00001100","11111011","00000101","11111000","11110001","11111011","00001000","11111000","11110011","11110010","11101111","11110101","00000101","11110011","11111101","11110001","00000001","00000101","11111001","11111000","00010000","11110010","00001011","00010000","11111111","00000010","11110011","00010000","00000000","11110101","11110101","00001000","00001011","11110010","00000100","00001001","11111001","11111110","11110110","11110111","11111000","00001101","11111011","00001000","00000100","11111101"),
        ("11111110","00000111","00010001","00010000","00011010","00000000","11110100","11111000","00000100","00001110","00000001","00001010","00001001","00000011","00001000","11111011","00001011","00000110","11111000","00000010","11111001","11110010","11110100","00000001","11110011","00001110","00001110","11101110","00000001","11100111","00000001","11111101","00000011","00010010","00010001","11111000","00000000","00001111","00000101","11111010","11111010","11111101","11111101","11101110","00000100","00011011","00011001","00001011","00001011","00001110","11111100","00001000","00000111","00010101","00001110","11110001","00000000","11110011","00001010","00010000","00000110","11110100","11111010","00000111"),
        ("00000110","00000000","00000010","00001100","11111011","11101100","11111000","00000011","00000101","11110100","00000000","00001100","00000010","00001100","00000011","00000101","00000110","11110100","00000101","00001100","11111111","11110100","11110011","11110101","00000100","00001110","00001011","11111001","00000100","11111110","11110101","11111010","11111100","00000010","00001101","11110010","11101111","00000010","00001100","00001110","00001001","11111000","00001110","11110000","11110110","00001011","11111100","11111101","00001001","11110101","00000011","00000010","11111100","11110110","11111110","00000111","11111011","11111111","00001010","11101111","11110100","11111100","00000100","00001010"),
        ("00000111","00000100","00001101","00011110","11111111","11111010","11111011","00001101","11111000","00001001","00000110","00000011","00011001","00011111","00000010","11110000","00000010","00010101","00011011","00011110","00011000","00101110","00010010","11110010","11110010","00001101","00011101","00010100","00001000","00001111","00000000","11110101","00001110","11110010","11111001","00000001","11101100","11110100","00001011","00000101","00001100","00001010","00000010","11111010","00000000","00000110","11110010","00000111","00000100","00000001","00011001","00010011","00001110","00010110","00001000","00001001","11111100","11110010","11101101","00000111","00101011","00001101","00000100","00010101")
    );
    constant WEIGHTS_2 : neural_matrix := (
        ("00000101","00000010","11111010","11101010","00100100","00001011","11111110","11111100","11111100","00010111","11111001","11111000","00000000","00001101","00001111","11110000","00001110","00001100","00001110","00011101"),
        ("00001100","00010111","00001010","00011101","11101011","00000010","11110100","11111001","00010110","00010001","00011001","11110111","11111111","00000010","11101010","00001101","00001011","11110011","00000100","00010111"),
        ("11111100","00000111","00010111","11101011","11110000","00001001","00010111","00000010","00000000","00010110","00011111","00001001","00000011","11110110","11111101","11100110","11111111","11111101","00000011","00001110"),
        ("11111111","11111001","11111100","00010001","11101011","00010100","00001000","00010011","11111011","11101100","00011010","00001111","00001000","11101110","00011100","11110010","11110011","00011001","00001001","11111110"),
        ("11111001","00000001","00000101","00001110","00100001","00000001","11111110","00000011","00010100","00011010","11110000","00001010","11110101","00010101","11100111","00010001","00001001","00000110","00001100","11110111"),
        ("00100101","00001011","11111001","00001100","00011010","00001001","00001111","11110010","11111101","11110010","00000010","00001111","00001000","11101100","11110101","00011000","00001001","00011010","00000010","11110111"),
        ("00001000","00000110","00100100","11101100","11110000","11111110","00001110","11111110","11111110","00011101","11110100","00001110","11111111","00010110","00001101","00011010","00001111","00001101","00001100","11111010"),
        ("00010001","00001000","11110111","00011010","11111110","00000011","00001100","00000000","00001111","11110101","11111110","00001001","11111101","00100110","00100110","11111101","11111001","11111110","11111101","11101000"),
        ("11110001","00010110","00001001","00010011","00001110","00000010","11110111","00000110","11110000","00001110","00001011","00001110","00000001","11110001","00010111","00010010","11110001","11111000","00000000","00010000"),
        ("11101110","11111101","11111000","00000011","00001010","00001110","00001110","00011111","00001111","11101010","11110110","11111110","00011000","00010100","00001101","00000111","00001100","11111011","00000110","00011101")
    );

    -- Enumerated structures of each weights-biases pair.
    -- NOTE: 'g_' prefix denotes "globality" in the Hungarian Notation.
    constant g_LAYER_1 : layer_parameters := (
        WEIGHTS_1,
        BIASES_1
    );
    constant g_LAYER_2 : layer_parameters := (
        WEIGHTS_2,
        BIASES_2
    );
    
    
    -- NOTE: There is no synth'able way to structure/group records,
    -- with variable-length elements, together in VHDL.  Unfortunately,
    -- dynamically allocated arrays, which would otherwise work here,
    -- are outright impossible to synthetize and nor can something like
    -- an "array of identifiers" help, either.
    -- A record of records could, technically, group these, but then
    -- again there is NO way to iterate over a record's elements.
    --
    -- The entire network comprising of the aforementioned layers
    --constant NETWORK_PARAMETERS : network_layers := 
    --    (g_LAYER_1, g_LAYER_2);
    
end package network_params;