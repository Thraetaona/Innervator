-- ---------------------------------------------------------------------
-- SPDX-License-Identifier: LGPL-3.0-or-later or CERN-OHL-W-2.0
-- uart_xmtr.vhd is a part of Innervator.
-- ---------------------------------------------------------------------


library ieee;
    use ieee.std_logic_1164.all;

library config;
    use config.constants.all;

-- TODO (when needed)
-- A simplex async. transmitter (in 8-N-1 frame)
architecture transmitter of uart is -- [RTL arch.]
    -- Placeholder
begin
    -- Placeholder
end architecture transmitter;


-- ---------------------------------------------------------------------
-- END OF FILE: uart_xmtr.vhd
-- ---------------------------------------------------------------------